// Vitis Shim requires no dynamically generated macros 
